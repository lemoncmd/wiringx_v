module wiringx

// init function for wiringx
fn init() {
}

// cleanup function for wiringx
fn cleanup() {
}
